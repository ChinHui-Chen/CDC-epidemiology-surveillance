BBC News | World | UK Edition$Sat, 11 Oct 2008 22:37:29 GMT
BBC News | News Front Page | UK Edition$Sat, 11 Oct 2008 22:37:29 GMT
CNN.com - Health$Fri, 10 Oct 2008 14:56:54 EDT

CNN.com - WORLD$Sat, 11 Oct 2008 19:19:34 EDT
CNN.com Recently Published/Updated$Sat, 11 Oct 2008 19:58:26 EDT
Google News - Top Stories$Sun, 12 Oct 2008 00:15:21 GMT
BBC News | Health | UK Edition$Sat, 11 Oct 2008 23:17:50 GMT
